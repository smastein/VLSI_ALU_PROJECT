module mtm_Alu_serializer (
    input wire clk,
	input wire rst_n,
	input wire C,
	input wire CTL_out,
	output reg sout
) ;

endmodule
